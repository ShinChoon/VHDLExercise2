

# LEF File for Accumulated Process Antenna Effects at the Boundary Pins
# *********************************************************************

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;

MACRO microcontroller_interface_8_8 
  PIN PC_tot[7] 
    ANTENNAPARTIALMETALAREA 1.2424 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.6196 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNAPARTIALMETALAREA 0.4584 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0916 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0162 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 46.4444 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 221.148 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 2.64198 LAYER Via5 ;
  END PC_tot[7]
  PIN PC_tot[6] 
    ANTENNAPARTIALMETALAREA 7.958 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 35.8398 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNAPARTIALMETALAREA 0.0264 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1476 LAYER Metal5 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via5 ;
    ANTENNAPARTIALMETALAREA 0.4512 LAYER Metal6 ;
    ANTENNAPARTIALMETALSIDEAREA 2.0592 LAYER Metal6 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0162 LAYER Metal6 ; 
    ANTENNAMAXAREACAR 82.1975 LAYER Metal6 ;
    ANTENNAMAXSIDEAREACAR 383.815 LAYER Metal6 ;
    ANTENNAMAXCUTCAR 2.94444 LAYER Via6 ;
  END PC_tot[6]
  PIN PC_tot[5] 
    ANTENNAPARTIALMETALAREA 8.0992 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 36.4752 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNAPARTIALMETALAREA 0.0528 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2952 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0162 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 75.5802 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 354.037 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 2.64198 LAYER Via5 ;
  END PC_tot[5]
  PIN PC_tot[4] 
    ANTENNAPARTIALMETALAREA 4.8044 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 21.6486 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02925 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 172.793 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 783.385 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 1.43932 LAYER Via4 ;
  END PC_tot[4]
  PIN PC_tot[3] 
    ANTENNAPARTIALMETALAREA 3.2764 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8014 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0162 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 218.469 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 995.259 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 2.33951 LAYER Via4 ;
  END PC_tot[3]
  PIN PC_tot[2] 
    ANTENNAPARTIALMETALAREA 7.0692 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 31.8402 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0162 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 457.136 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 2067.48 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 2.33951 LAYER Via4 ;
  END PC_tot[2]
  PIN PC_tot[1] 
    ANTENNAPARTIALMETALAREA 6.9364 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 31.2426 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02925 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 245.737 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 1111.63 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 1.43932 LAYER Via4 ;
  END PC_tot[1]
  PIN PC_tot[0] 
    ANTENNAPARTIALMETALAREA 11.0992 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 50.004 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.07785 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 162.168 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 737.017 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 2.89198 LAYER Via4 ;
  END PC_tot[0]
  PIN instruction_in[13] 
    ANTENNAPARTIALMETALAREA 1.9556 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 8.829 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02925 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 69.2274 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 316.133 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.3094 LAYER Via3 ;
  END instruction_in[13]
  PIN instruction_in[12] 
    ANTENNAPARTIALMETALAREA 3.4804 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6906 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02925 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 121.32 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 550.769 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.27179 LAYER Via3 ;
  END instruction_in[12]
  PIN instruction_in[11] 
    ANTENNAPARTIALMETALAREA 1.702 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6878 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02925 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 60.5197 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 277.169 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.27179 LAYER Via3 ;
  END instruction_in[11]
  PIN instruction_in[10] 
    ANTENNAPARTIALMETALAREA 2.1948 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 9.9054 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02925 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 76.694 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 349.733 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.3094 LAYER Via3 ;
  END instruction_in[10]
  PIN instruction_in[9] 
    ANTENNAPARTIALMETALAREA 2.5956 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.7378 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0909 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 43.0082 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 200.203 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAMAXCUTCAR 3.50761 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 1.8192 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 8.2152 LAYER Metal4 ;
    ANTENNAGATEAREA 0.16875 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 53.7886 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 248.885 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 6.57716 LAYER Via4 ;
  END instruction_in[9]
  PIN instruction_in[8] 
    ANTENNAPARTIALMETALAREA 1.7004 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6806 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02925 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 62.5812 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 286.226 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.3094 LAYER Via3 ;
  END instruction_in[8]
  PIN instruction_in[7] 
    ANTENNAPARTIALMETALAREA 2.9604 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.3218 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0098 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 1.1152 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.076 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0747 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 36.5375 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 174.212 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 9.45328 LAYER Via4 ;
  END instruction_in[7]
  PIN instruction_in[6] 
    ANTENNAPARTIALMETALAREA 2.6164 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 11.8026 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02925 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 96.0034 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 436.626 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.3094 LAYER Via3 ;
  END instruction_in[6]
  PIN instruction_in[5] 
    ANTENNAPARTIALMETALAREA 2.3828 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7514 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02925 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 83.1214 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 378.656 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.3094 LAYER Via3 ;
  END instruction_in[5]
  PIN instruction_in[4] 
    ANTENNAPARTIALMETALAREA 3.4184 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 15.4116 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02925 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 126.048 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 571.826 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 1.3094 LAYER Via3 ;
  END instruction_in[4]
  PIN instruction_in[3] 
    ANTENNAPARTIALMETALAREA 3.9392 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.8416 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.12645 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 70.9022 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 327.8 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAMAXCUTCAR 7.5583 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 1.4088 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.3684 LAYER Metal4 ;
    ANTENNAGATEAREA 0.22365 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 77.2014 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 356.275 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 7.5583 LAYER Via4 ;
  END instruction_in[3]
  PIN instruction_in[2] 
    ANTENNAPARTIALMETALAREA 4.804 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 21.762 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 72.3887 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 333.324 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 4.94444 LAYER Via3 ;
  END instruction_in[2]
  PIN instruction_in[1] 
    ANTENNAPARTIALMETALAREA 4.1564 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 18.7902 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1881 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 81.9126 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 378.006 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 9.84259 LAYER Via3 ;
  END instruction_in[1]
  PIN instruction_in[0] 
    ANTENNAPARTIALMETALAREA 2.3472 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5624 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 1.0288 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.6584 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04545 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 47.3768 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 221.43 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 4.5183 LAYER Via4 ;
  END instruction_in[0]
  PIN opcode_status[1] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 4.5264 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 20.3976 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2367 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 41.4069 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 193.99 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END opcode_status[1]
  PIN opcode_status[0] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 4.398 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8198 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2367 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 32.0032 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 182.573 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.3159 LAYER Via4 ;
  END opcode_status[0]
  PIN statusOutSPI[2] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.1024 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4896 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 13.2435 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 98.1551 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END statusOutSPI[2]
  PIN statusOutSPI[1] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.0312 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1404 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 22.4068 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 139.39 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2531 LAYER Via4 ;
  END statusOutSPI[1]
  PIN statusOutSPI[0] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.0312 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.1404 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 23.8776 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 146.008 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END statusOutSPI[0]
  PIN resultOutMemSPI[7] 
    ANTENNAPARTIALMETALAREA 2.9072 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 13.0824 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.1928 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8964 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 4.4104 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.8756 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 32.8753 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 186.629 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2875 LAYER Via5 ;
  END resultOutMemSPI[7]
  PIN resultOutMemSPI[6] 
    ANTENNADIFFAREA 2.62222 LAYER Metal3 ; 
    ANTENNAPARTIALMETALAREA 7.3296 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 33.012 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 45.6122 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 243.684 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 12.2308 LAYER Via3 ;
  END resultOutMemSPI[6]
  PIN resultOutMemSPI[5] 
    ANTENNAPARTIALMETALAREA 3.2936 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 14.8212 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.1776 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.828 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 3.4824 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6996 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 32.9501 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 186.966 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2753 LAYER Via5 ;
  END resultOutMemSPI[5]
  PIN resultOutMemSPI[4] 
    ANTENNAPARTIALMETALAREA 2.3968 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 10.7856 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.0864 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4176 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 4.6984 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 21.1716 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 42.878 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 231.641 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2875 LAYER Via5 ;
  END resultOutMemSPI[4]
  PIN resultOutMemSPI[3] 
    ANTENNAPARTIALMETALAREA 3.7736 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 16.9812 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.1928 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.8964 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 3.3536 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 15.12 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 40.4748 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 220.827 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2753 LAYER Via5 ;
  END resultOutMemSPI[3]
  PIN resultOutMemSPI[2] 
    ANTENNAPARTIALMETALAREA 1.7056 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.6752 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.0864 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.4176 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 4.5384 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 20.4516 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 54.8617 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 285.567 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2875 LAYER Via5 ;
  END resultOutMemSPI[2]
  PIN resultOutMemSPI[1] 
    ANTENNAPARTIALMETALAREA 1.6352 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.3584 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 1.3176 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.958 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 5.8504 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 26.3556 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 53.507 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 279.472 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2753 LAYER Via5 ;
  END resultOutMemSPI[1]
  PIN resultOutMemSPI[0] 
    ANTENNAPARTIALMETALAREA 1.7568 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9056 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 5.1656 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 23.274 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 5.3224 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 23.9796 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 38.922 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 213.839 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2753 LAYER Via5 ;
  END resultOutMemSPI[0]
  PIN addrSPI[7] 
    ANTENNADIFFAREA 0.1448 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.0464 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.2088 LAYER Metal4 ;
  END addrSPI[7]
  PIN addrSPI[6] 
    ANTENNADIFFAREA 3.57945 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 18.722 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 84.249 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.285975 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 81.2253 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 404.064 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 11.8622 LAYER Via4 ;
  END addrSPI[6]
  PIN addrSPI[5] 
    ANTENNADIFFAREA 3.57945 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 19.0296 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 85.662 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.285975 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 80.4238 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 400.556 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 11.865 LAYER Via4 ;
  END addrSPI[5]
  PIN addrSPI[4] 
    ANTENNADIFFAREA 0.572 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 14.6252 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 65.871 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0585 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 270.166 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 1248.89 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 9.2547 LAYER Via4 ;
  END addrSPI[4]
  PIN addrSPI[3] 
    ANTENNADIFFAREA 3.57945 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 19.344 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 87.0768 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.285975 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 83.5262 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 414.519 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 11.8622 LAYER Via4 ;
  END addrSPI[3]
  PIN addrSPI[2] 
    ANTENNADIFFAREA 3.57945 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 19.396 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 87.3108 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.285975 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 83.5542 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 414.643 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 11.865 LAYER Via4 ;
  END addrSPI[2]
  PIN addrSPI[1] 
    ANTENNAPARTIALMETALAREA 16.9052 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 76.0734 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNADIFFAREA 3.57945 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 4.2336 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 19.08 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.285975 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 37.3291 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 206.731 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 11.8822 LAYER Via5 ;
  END addrSPI[1]
  PIN addrSPI[0] 
    ANTENNAPARTIALMETALAREA 17.152 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 77.2128 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNADIFFAREA 3.57945 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 5.0824 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 22.8996 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.285975 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 37.4075 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 207.083 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 11.8822 LAYER Via5 ;
  END addrSPI[0]
  PIN Instruction[4] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.3384 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.0228 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 56.776 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 293.921 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2531 LAYER Via4 ;
  END Instruction[4]
  PIN Instruction[3] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.3336 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 6.03 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 23.6454 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 144.963 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END Instruction[3]
  PIN Instruction[2] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.8976 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 4.0392 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 24.4871 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 148.751 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END Instruction[2]
  PIN Instruction[1] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.1408 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 5.1336 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 65.9805 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 335.341 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2531 LAYER Via4 ;
  END Instruction[1]
  PIN Instruction[0] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 0.3456 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 1.584 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 16.868 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 114.465 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END Instruction[0]
  PIN PC_out[7] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.4824 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.6708 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 52.5746 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 275.015 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2531 LAYER Via4 ;
  END PC_out[7]
  PIN PC_out[6] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.4056 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.3252 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 51.2082 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 268.865 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END PC_out[6]
  PIN PC_out[5] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.2696 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.7132 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 49.8136 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 262.59 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2531 LAYER Via4 ;
  END PC_out[5]
  PIN PC_out[4] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.7824 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.5208 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 49.0807 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 259.293 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2531 LAYER Via4 ;
  END PC_out[4]
  PIN PC_out[3] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.1632 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.2344 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 45.5483 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 243.396 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END PC_out[3]
  PIN PC_out[2] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.8432 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.7944 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 41.434 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 224.882 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END PC_out[2]
  PIN PC_out[1] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.7064 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.1788 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 38.044 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 209.627 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2531 LAYER Via4 ;
  END PC_out[1]
  PIN PC_out[0] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.4784 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.1528 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 34.2612 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 192.604 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END PC_out[0]
  PIN A_out[7] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.3424 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.5408 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 34.2794 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 192.686 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END A_out[7]
  PIN A_out[6] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.2656 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 10.1952 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 33.4304 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 188.865 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END A_out[6]
  PIN A_out[5] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.1904 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.8568 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 31.3537 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 179.521 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2531 LAYER Via4 ;
  END A_out[5]
  PIN A_out[4] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.0528 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.2376 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 27.6689 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 162.939 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END A_out[4]
  PIN A_out[3] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.6728 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.5276 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 26.7546 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 158.824 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END A_out[3]
  PIN A_out[2] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.7732 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9794 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 24.7088 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 149.619 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2531 LAYER Via4 ;
  END A_out[2]
  PIN A_out[1] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.0924 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 9.4158 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 23.0848 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 142.31 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2653 LAYER Via4 ;
  END A_out[1]
  PIN A_out[0] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 1.7588 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 7.9146 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2205 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 21.3347 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 134.435 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2531 LAYER Via4 ;
  END A_out[0]
  PIN W_out[7] 
    ANTENNAPARTIALMETALAREA 2.6416 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.916 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.14265 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 58.8725 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 275.737 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0098 LAYER Via4 ;
    ANTENNAMAXCUTCAR 4.91181 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 1.7632 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.992 LAYER Metal5 ;
    ANTENNAGATEAREA 0.4086 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 63.1877 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 295.296 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2875 LAYER Via5 ;
  END W_out[7]
  PIN W_out[6] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 2.656 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 11.9808 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.40545 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 33.8174 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 182.128 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.3329 LAYER Via4 ;
  END W_out[6]
  PIN W_out[5] 
    ANTENNAPARTIALMETALAREA 2.8688 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 12.9384 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.04545 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 101.303 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 467.203 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNAMAXCUTCAR 3.2617 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 0.3784 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 1.7316 LAYER Metal5 ;
    ANTENNAGATEAREA 0.31455 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 102.506 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 472.708 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2847 LAYER Via5 ;
  END W_out[5]
  PIN W_out[4] 
    ANTENNAPARTIALMETALAREA 3.3852 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 15.2334 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 1.7208 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 7.7724 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.3699 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 21.8503 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 136.963 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2875 LAYER Via5 ;
  END W_out[4]
  PIN W_out[3] 
    ANTENNAPARTIALMETALAREA 3.5744 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 16.0848 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0162 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 236.395 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 1077.52 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNAMAXCUTCAR 3.92593 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 1.0648 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 4.8204 LAYER Metal5 ;
    ANTENNAGATEAREA 0.35685 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 239.379 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1091.03 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2789 LAYER Via5 ;
  END W_out[3]
  PIN W_out[2] 
    ANTENNAPARTIALMETALAREA 3.2392 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 14.5764 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNADIFFAREA 2.62222 LAYER Metal5 ; 
    ANTENNAPARTIALMETALAREA 1.1768 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 5.3244 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.28215 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 24.3606 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 127.77 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 12.2696 LAYER Via5 ;
  END W_out[2]
  PIN W_out[1] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 4.1472 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 18.6912 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.37305 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 28.6546 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 167.412 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2462 LAYER Via4 ;
  END W_out[1]
  PIN W_out[0] 
    ANTENNADIFFAREA 2.62222 LAYER Metal4 ; 
    ANTENNAPARTIALMETALAREA 3.816 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 17.172 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2952 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 36.1678 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 169.533 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 12.2531 LAYER Via4 ;
  END W_out[0]
  PIN clk 
    ANTENNAPARTIALMETALAREA 0.0092 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 0.0414 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.0788 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.3834 LAYER Metal4 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.08775 LAYER Metal4 ; 
    ANTENNAMAXAREACAR 17.2274 LAYER Metal4 ;
    ANTENNAMAXSIDEAREACAR 80.3795 LAYER Metal4 ;
    ANTENNAMAXCUTCAR 0.651852 LAYER Via4 ;
  END clk
  PIN rst 
    ANTENNAPARTIALMETALAREA 1.322 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 5.9778 LAYER Metal3 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.0162 LAYER Metal3 ; 
    ANTENNAMAXAREACAR 86.7716 LAYER Metal3 ;
    ANTENNAMAXSIDEAREACAR 404.148 LAYER Metal3 ;
    ANTENNAMAXCUTCAR 3.25309 LAYER Via3 ;
  END rst
  PIN instr_wr 
    ANTENNAPARTIALMETALAREA 3.8384 LAYER Metal3 ;
    ANTENNAPARTIALMETALSIDEAREA 17.2728 LAYER Metal3 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via3 ;
    ANTENNAPARTIALMETALAREA 0.1472 LAYER Metal4 ;
    ANTENNAPARTIALMETALSIDEAREA 0.6912 LAYER Metal4 ;
    ANTENNAPARTIALCUTAREA 0.0049 LAYER Via4 ;
    ANTENNAPARTIALMETALAREA 6.5384 LAYER Metal5 ;
    ANTENNAPARTIALMETALSIDEAREA 29.4516 LAYER Metal5 ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.02925 LAYER Metal5 ; 
    ANTENNAMAXAREACAR 236.68 LAYER Metal5 ;
    ANTENNAMAXSIDEAREACAR 1071.64 LAYER Metal5 ;
    ANTENNAMAXCUTCAR 1.64444 LAYER Via5 ;
  END instr_wr
END microcontroller_interface_8_8

END LIBRARY
