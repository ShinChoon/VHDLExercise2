/prog/cadence/gpdk/g045/GPDK045/gsclib045_all_v4.4/gsclib045_tech/lef/gsclib045_tech.lef