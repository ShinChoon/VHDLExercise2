/prog/cadence/gpdk/g045/GPDK045/gsclib045_all_v4.4/gsclib045_lvt/lef/gsclib045_lvt_macro.lef